library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;


entity vga_sync is
	port(
		clk, reset : in std_logic;
		hsync, vsync : out std_logic;
		video_on, p_tick : out std_logic;
		pixel_x, pixel_y : out std_logic_vector(9 downto 0)
		);
		
end vga_sync;

architecture arch of vga_sync is

	constant HD : integer := 640; --horizontal display area 640
	constant HF : integer := 16; --				 front porch 16
	constant HB : integer := 48; --			  	 back porch 48
	constant HR : integer := 96;	--           retrace 96
	
	constant VD : integer := 480; --vertical display area 480
	constant VF : integer := 10; --		  	  front porch 10
	constant VB : integer := 33; --		 	  back porch 33
	constant VR : integer := 2; --           retrace 2

	signal mod2_reg, mod2_next : std_logic;
	
	signal v_count_reg, v_count_next : unsigned(9 downto 0);
	signal h_count_reg, h_count_next : unsigned(9 downto 0);
	
	signal v_sync_reg, v_sync_next : std_logic;
	signal h_sync_reg, h_sync_next : std_logic;
	
	signal h_end, v_end, pixel_tick : std_logic;


begin
	
	process(clk, reset)
	begin
		
		if (reset='1') then
		 	mod2_reg <= '0';
			v_count_reg <= (others => '0');
			h_count_reg <= (others => '0');
			v_sync_reg <= '0';
			h_sync_reg <= '0';
		elsif (rising_edge(clk)) then
			mod2_reg <= mod2_next;
			v_count_reg <= v_count_next;
			h_count_reg <= h_count_next;
			v_sync_reg <= v_sync_next;
			h_sync_reg <= h_sync_next;
		end if;
		
	end process;
	
	mod2_next <= not(mod2_reg);
	pixel_tick <= '1' when mod2_reg = '1' else '0';
	
	h_end <= '1' when h_count_reg = (HD + HF + HB + HR -1) else '0';
	v_end <= '1' when v_count_reg = (VD + VF + VB + VR -1) else '0';
	
	process (h_count_reg, h_end, pixel_tick)
	begin
		if (pixel_tick = '1') then
			if (h_end = '1') then
				h_count_next <= (others => '0');
			else
				h_count_next <= h_count_reg +1;
			end if;
		else
			h_count_next <= h_count_reg ;
		end if;
	end process;
	
	process (v_count_reg, v_end, pixel_tick, h_end)
	begin
		if (pixel_tick = '1' and h_end ='1') then
			if (v_end = '1') then
				v_count_next <= (others => '0');
			else
				v_count_next <= v_count_reg +1;
			end if;
		else
			v_count_next <= v_count_reg ;
		end if;
	end process;
	
	h_sync_next <=
		'1' when ((h_count_reg >= (HD + HF)) and (h_count_reg <= (HD + HF + HR -1))) else    --(h_count_reg >= (HD + HF)) and (h_count_reg <= (HD + HF + HR -1))
		'0';
	
	v_sync_next <=
		'1' when ((v_count_reg >= (VD + VF)) and (v_count_reg <= (VD + VF + VR -1))) else    --(v_count_reg >= (VD + VF)) and (v_count_reg <= (VD + VF + VR -1))
		'0';
		
	video_on <=
		'1' when ((h_count_reg < HD) and (v_count_reg < VD)) else
		'0';
		
	hsync <= h_sync_reg;
	vsync <= v_sync_reg;
	pixel_x <= std_logic_vector(h_count_reg);
	pixel_y <= std_logic_vector(v_count_reg);
	p_tick <= pixel_tick;
	
	
end arch;

